module andgate(a,b,y);
input a;
input b;
output y;
reg y;

and a1(y,a,b);

endmodule
