class and_transaction;
//PROPERTIES
//INPUTS declare as rand variables
  rand bit [1:0] a;
  rand bit [1:0] b;
  //Output
  bit y;
